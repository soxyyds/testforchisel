module nihao ();
helloworld
#(
    .WIDTH(8)
) dut (
    .in1(in1),
    .in2(in2),
    .out(out)
);
endmodule

//更新一次
