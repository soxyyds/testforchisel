module test ();

endmodule
